﻿return {

help_title = "cmd_pm2offliners.lua",
help_usage = "[+!#]pm add <ANVÄNDARNAMN> <MEDDELANDE>  / eller: [+!#]pm del",
help_desc = "Skickar ett PM till en frånkopplad registrerad användare",

ucmd_menu_add_1 = "Användare",
ucmd_menu_add_2 = "Meddelande",
ucmd_menu_add_3 = "PM till Frånkopplad",
ucmd_menu_add_4 = "skicka meddelande",
ucmd_menu_add_5 = "till ANVÄNDARNAMN från lista",
ucmd_menu_add_6 = { "Användare", "Meddelande", "PM till Frånkopplad", "skicka meddelande", "till ANVÄNDARNAMN" },
ucmd_menu_del = { "Användare", "Meddelande", "PM till Frånkopplad", "ta bort databas" },
ucmd_popup = "Meddelande:",
ucmd_popup2 = "Användarnamn:",

msg_denied = "Du har inte behörighet att använda detta kommando.",
msg_usage = "Användning: [+!#]pm add <ANVÄNDARNAMN> <MEDDELANDE>  / eller: [+!#]pm del",
msg_fail_1 = "Användaren är inte registrerad.",
msg_fail_2 = "Användaren är redan ansluten.",
msg_ok = "Meddelandet är sparat.",
msg_del_1 = "Databasen har rensats.",
msg_del_2 = "Databasen är redan tom.",
msg_reply = "Du har fått [%s] meddelande(n) medans du var frånkopplad.",
msg_pm_1 = "Frånkopplade PM %s  |  ",
msg_pm_2 = "Avsändare: %s  |  Datum: %s \n\n",
msg_pm_3 = "Meddelande: %s \n\n",
msg_confirm = "Det privata meddelandet du skickade till  %s  har mottagits.\n\nDatum: %s\nMeddelande: %s",

}
return {

    msg_too_many_slots = "Du har för många slottar öppnade. En användare med %s får ha maximalt %s slottar öppnade. Du hade %s slottar.",
    msg_too_few_slots = "Du har för få slottar öppnade. En användare med %s måste ha minst %s slottar öppnade. Du hade %s slottar.",
    msg_too_many_hubs = "Du är i för många hubbar. En användare med %s får vara ansluten till maximalt %s hubbar samtidigt. Du var ansluten till %s hubbar.",

    msg_ban = "%s har blivit bannad och kickad av %s i %s minuter därför att: %s",

}

return {

    help_title = "Banner",
    help_usage = "[+!#]banner [show|set_msg <text>|set_time <tid>]",
    help_desc = "[show] visar bannern | [set_msg <text>] ange <text> som bannertext | [set_time <tid>] ange <tid> som tidsinterval.",

    msg_denied = "Du har inte behörighet att använda detta kommando.",
    msg_usage = "Användning: [+!#]banner show och [+!#]banner set_msg <text> och [+!#]banner set_time <tid>",
    msg_time = "Bannern skickas ut var %s timme.",

    ucmd_menu_show = { "Hubb", "etc", "Banner", "Visa Banner" },
    ucmd_menu_set_msg = { "Hubb", "etc", "Banner", "Ange Banner" },
    ucmd_menu_set_time = { "Hubb", "etc", "Banner", "Ange Intervall" },

    ucmd_popup1 = "Ange den nya texten.",
    ucmd_popup2 = "Ange tidsintervallen (i timmar).",

}